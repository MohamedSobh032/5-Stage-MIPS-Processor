LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY ControlUnit IS
	PORT (
		---------------- INSTRUCTION OPCODE ----------------
		INSTRUCTION : IN STD_LOGIC_VECTOR(4 DOWNTO 0);

		---------------- CONTROL SIGNALS ----------------
		-- WRITE BACK 1 		--> 0
		-- WRITE BACK 2 		--> 1
		-- Z/N F			--> 2
		-- C/OV F       		--> 3
		-- MemRead			--> 4
		-- MemWrite			--> 5
		-- FREE				--> 6
		-- PROTECT			--> 7
		-- IMMEDIATE    		--> 8
		-- BRANCH			--> 9
		-- BRANCH ZERO 			--> 10
		-- SP DEC 			--> 11
		-- SP INC 			--> 12
		-- OUTPUT PORT  		--> 13
		-- INPUT PORT   		--> 14
		-- STORE        		--> 15
		-- PC SAVE/GET  		--> 16
		-- LENGTH EXT   		--> 17
		-- First Operand Dependency 	--> 18
		-- Second Operand Dependency	--> 19
		-- Push the CCR			--> 20
		-- Pop the PC			--> 21
		CONTROL_SIGNALS : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);

		---------------- ALU OPCODE ----------------
		-- NOT  --> 0001
		-- NEG  --> 0010
		-- INC  --> 0011
		-- DEC  --> 0100
		-- ADD  --> 0101
		-- ADDI --> 0101
		-- SUB  --> 0110
		-- SUBI --> 0110
		-- AND  --> 0111
		-- OR   --> 1000
		-- XOR  --> 1001
		-- CMP  --> 1010
		-- LDM  --> 1011
		-- LDD  --> 0101
		-- STD  --> 0101
		ALU_OPCODE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE a_ControlUnit OF ControlUnit IS
	BEGIN
		---- ALU OPCODE SIGNAL SELECTION ----
		WITH INSTRUCTION SELECT
			ALU_OPCODE <=
				"0001" WHEN "00001", -- NOT
				"0010" WHEN "00010", -- NEG
				"0011" WHEN "00011", -- INC
				"0100" WHEN "00100", -- DEC
				"0101" WHEN "01001", -- ADD
				"0101" WHEN "01010", -- ADDI
				"0110" WHEN "01011", -- SUB
				"0110" WHEN "01100", -- SUBI
				"0111" WHEN "01101", -- AND
				"1000" WHEN "01110", -- OR
				"1001" WHEN "01111", -- XOR
				"0110" WHEN "10000", -- CMP
				"1011" WHEN "10011", -- LDM
				"0101" WHEN "10100", -- LDD
				"0101" WHEN "10101", -- STD
				"0000" WHEN OTHERS;
		
		---- CONTROL SIGNAL SELECTION ----
		WITH INSTRUCTION SELECT
			CONTROL_SIGNALS <=
				"000000000000000000000000" WHEN "00000",	-- NOP
				"000001000000000000000101" WHEN "00001",	-- NOT
				"000001000000000000001101" WHEN "00010",	-- NEG
				"000001000000000000001101" WHEN "00011",	-- INC
				"000001000000000000001101" WHEN "00100",	-- DEC
				"000001000010000000000000" WHEN "00101",	-- OUT
				"000000000100000000000001" WHEN "00110",	-- IN
				"000001000000000000000001" WHEN "00111",	-- MOV
				"000011000000000000000011" WHEN "01000",	-- SWAP
				"000011000000000000001101" WHEN "01001",	-- ADD
				"000001000000000100001101" WHEN "01010",	-- ADDI
				"000011000000000000001101" WHEN "01011",	-- SUB
				"000001000000000100001101" WHEN "01100",	-- SUBI
				"000011000000000000000101" WHEN "01101",	-- AND
				"000011000000000000000101" WHEN "01110",	-- OR
				"000011000000000000000101" WHEN "01111",	-- XOR
				"000011000000000000000100" WHEN "10000",	-- CMP
				"000001000000100000100000" WHEN "10001",	-- PUSH
				"000000000001000000010001" WHEN "10010",	-- POP
				"000000100000000100000001" WHEN "10011",	-- LDM
				"000011000000000100010001" WHEN "10100",	-- LDD
				"000011001000000100100000" WHEN "10101",	-- STD
				"000000000000000010000000" WHEN "10110",	-- PROT
				"000000000000000001000000" WHEN "10111",	-- FREE
				"000001000000010000000000" WHEN "11000",	-- JZ
				"000001000000001000000000" WHEN "11001",	-- JMP
				"000001010000101000100000" WHEN "11010",	-- CALL
				"101000010001000000010000" WHEN "11011",	-- RET
				"000000010001001000010000" WHEN "11100",	-- RTI
				"000100010000100000100000" WHEN "11101",	-- INT_PC
				"001000010000100000101100" WHEN "11110",	-- INT_CCR
				"010000000001000000011100" WHEN "11111",	-- POP_CCR
				(OTHERS => '0') WHEN OTHERS;

END a_ControlUnit;