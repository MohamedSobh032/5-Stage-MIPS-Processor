LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MemUseUnit IS
	PORT (
		-- CURRENT ADDRESSES IN THE EXECUTE --
		Rsrc1Addr     : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Rsrc2Addr     : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		-- ADDRESSES PERVIOUSLY IN EXECUTION STAGE --
		Rdst1Addr_MEM : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		MEM_READ      : IN STD_LOGIC;
		-- DEPENDENCY
		FIRST_DEPENDENCY  : IN STD_LOGIC;
		SECOND_DEPENDENCY : IN STD_LOGIC;
		-- STALL SIGNAL
		STALL         : OUT STD_LOGIC
	);
END MemUseUnit;


ARCHITECTURE a_MemUseUnit OF MemUseUnit IS

	SIGNAL COND_FIRST_OP  : STD_LOGIC;
	SIGNAL COND_SECOND_OP : STD_LOGIC;

	BEGIN
		COND_FIRST_OP  <= '1' WHEN ((Rsrc1Addr = Rdst1Addr_MEM) AND (MEM_READ = '1') AND (FIRST_DEPENDENCY  = '1')) ELSE '0';
		COND_SECOND_OP <= '1' WHEN ((Rsrc2Addr = Rdst1Addr_MEM) AND (MEM_READ = '1') AND (SECOND_DEPENDENCY = '1')) ELSE '0';
		STALL          <= '1' WHEN ((COND_FIRST_OP = '1') OR (COND_SECOND_OP = '1')) ELSE '0';

END ARCHITECTURE;

