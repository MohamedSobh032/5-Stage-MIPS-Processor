LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY ControlUnit IS
	PORT (
		---------------- INSTRUCTION OPCODE ----------------
		INSTRUCTION : IN STD_LOGIC_VECTOR(4 DOWNTO 0);

		---------------- CONTROL SIGNALS ----------------
		-- WRITE BACK 1 --> 0
		-- WRITE BACK 2 --> 1
		-- Z/N F	--> 2
		-- C/OV F       --> 3
		-- MemRead	--> 4
		-- MemWrite	--> 5
		-- FREE		--> 6
		-- PROTECT	--> 7
		-- IMMEDIATE    --> 8
		-- BRANCH	--> 9
		-- BRANCH ZERO 	--> 10
		-- SP OPERATION --> 11
		-- OUTPUT PORT  --> 12
		-- INPUT PORT   --> 13
		-- STORE        --> 14
		-- PC SAVE/GET  --> 15
		-- LENGTH EXT   --> 16
		CONTROL_SIGNALS : OUT STD_LOGIC_VECTOR(16 DOWNTO 0);

		---------------- ALU OPCODE ----------------
		-- NOT  --> 0001
		-- NEG  --> 0010
		-- INC  --> 0011
		-- DEC  --> 0100
		-- ADD  --> 0101
		-- ADDI --> 0101
		-- SUB  --> 0110
		-- SUBI --> 0110
		-- AND  --> 0111
		-- OR   --> 1000
		-- XOR  --> 1001
		-- CMP  --> 1010
		-- LDM  --> 1011
		-- LDD  --> 0101
		-- STD  --> 0101
		ALU_OPCODE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE a_ControlUnit OF ControlUnit IS
	BEGIN
		---- ALU OPCODE SIGNAL SELECTION ----
		WITH INSTRUCTION SELECT
			ALU_OPCODE <=
				"0001" WHEN "00001", -- NOT
				"0010" WHEN "00010", -- NEG
				"0011" WHEN "00011", -- INC
				"0100" WHEN "00100", -- DEC
				"0101" WHEN "01001", -- ADD
				"0101" WHEN "01010", -- ADDI
				"0110" WHEN "01011", -- SUB
				"0110" WHEN "01100", -- SUBI
				"0111" WHEN "01101", -- AND
				"1000" WHEN "01110", -- OR
				"1001" WHEN "01111", -- XOR
				"0110" WHEN "10000", -- CMP
				"1011" WHEN "10011", -- LDM
				"0101" WHEN "10100", -- LDD
				"0101" WHEN "10101", -- STD
				"0000" WHEN OTHERS;
		
		---- CONTROL SIGNAL SELECTION ----
		WITH INSTRUCTION SELECT
			CONTROL_SIGNALS <=
				"00000000000000000" WHEN "00000",	-- NOP
				"00000000000000101" WHEN "00001",	-- NOT
				"00000000000001101" WHEN "00010",	-- NEG
				"00000000000001101" WHEN "00011",	-- INC
				"00000000000001101" WHEN "00100",	-- DEC
				"00001000000000000" WHEN "00101",	-- OUT
				"00010000000000001" WHEN "00110",	-- IN
				"00000000000000001" WHEN "00111",	-- MOV
				"00000000000000011" WHEN "01000",	-- SWAP
				"00000000000001101" WHEN "01001",	-- ADD
				"00000000100001101" WHEN "01010",	-- ADDI
				"00000000000001101" WHEN "01011",	-- SUB
				"00000000100001101" WHEN "01100",	-- SUBI
				"00000000000000101" WHEN "01101",	-- AND
				"00000000000000101" WHEN "01110",	-- OR
				"00000000000000101" WHEN "01111",	-- XOR
				"00000000000000100" WHEN "10000",	-- CMP
				"00000100000100000" WHEN "10001",	-- PUSH
				"00000100000010001" WHEN "10010",	-- POP
				"10000000100000001" WHEN "10011",	-- LDM
				"00000000100010001" WHEN "10100",	-- LDD
				"00100000100100000" WHEN "10101",	-- STD
				"00000000010000000" WHEN "10110",	-- PROTECT
				"00000000001000000" WHEN "10111",	-- FREE
				"00000010000000000" WHEN "11000",	-- JZ
				"00000001000000000" WHEN "11001",	-- JMP
				"01000101000100000" WHEN "11010",	-- CALL
				"01000101000010000" WHEN "11011",	-- RET
				"01000101000010000" WHEN "11100",	-- RTI
				(OTHERS => '0') WHEN OTHERS;

END a_ControlUnit;