LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY OurALU IS
	PORT (
		CLK    : IN  STD_LOGIC;

		OpCode : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		
		Rsrc1  : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Rsrc2  : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Rdst   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		-- (3 = OVF) (2 = CF) (1 = NF) (0 = ZF)
		CCR    : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END OurALU;

ARCHITECTURE a_OurALU OF OurALU IS

	-------------------- MAIN COMPONENTS --------------------
	COMPONENT ALU_not IS
		PORT (
			Rsrc : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Rdst : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			Carry : OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT ALU_dec IS
		PORT (
			Rsrc : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Rdst : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			Carry : OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT ALU_or IS
		PORT (
			Rsrc1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Rsrc2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Rdst  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			Carry : OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT ALU_ldm IS
		PORT (
			Rsrc : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Rdst : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			Carry : OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT ALU_mov IS
		PORT (
			Rsrc : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Rdst : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			Carry : OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT ALU_cmp IS
		PORT (
			Rsrc1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Rsrc2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Rdst  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			Carry : OUT STD_LOGIC
		);
	END COMPONENT;

	-- OUTPUTS
	SIGNAL ALU_NOT_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ALU_DEC_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ALU_OR_OUT  : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ALU_LDM_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ALU_MOV_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ALU_CMP_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);

	-- CARRIES
	SIGNAL ALU_NOT_CARRY : STD_LOGIC;
	SIGNAL ALU_DEC_CARRY : STD_LOGIC;
	SIGNAL ALU_OR_CARRY  : STD_LOGIC;
	SIGNAL ALU_LDM_CARRY : STD_LOGIC;
	SIGNAL ALU_MOV_CARRY : STD_LOGIC;
	SIGNAL ALU_CMP_CARRY : STD_LOGIC;

	SIGNAL Mout : STD_LOGIC_VECTOR(31 DOWNTO 0);

	BEGIN

		u1  : ALU_not PORT MAP(Rsrc1,        ALU_NOT_OUT, ALU_NOT_CARRY);
		u4  : ALU_dec PORT MAP(Rsrc1,        ALU_DEC_OUT, ALU_DEC_CARRY);
		u7  : ALU_mov PORT MAP(Rsrc1,        ALU_MOV_OUT, ALU_MOV_CARRY);
		u14 : ALU_or  PORT MAP(Rsrc1, Rsrc2, ALU_OR_OUT , ALU_OR_CARRY);
		u16 : ALU_cmp PORT MAP(Rsrc1, Rsrc2, ALU_CMP_OUT, ALU_CMP_CARRY);
		u19 : ALU_ldm PORT MAP(Rsrc1,        ALU_LDM_OUT, ALU_LDM_CARRY);

		PROCESS (CLK)
		BEGIN
			IF rising_edge(CLK) THEN
				-- OUTPUT AND CARRY
				CASE OpCode IS
					WHEN "00001" =>
						Mout   <= ALU_NOT_OUT;
						CCR(2) <= ALU_NOT_CARRY;

					WHEN "00100" =>
						Mout   <= ALU_DEC_OUT;
						CCR(2) <= ALU_DEC_CARRY;

					WHEN "00111" =>
						Mout   <= ALU_MOV_OUT;
						CCR(2) <= ALU_MOV_CARRY;

					WHEN "01110" =>
						Mout   <= ALU_OR_OUT;
						CCR(2) <= ALU_OR_CARRY;
				
					WHEN "10000" =>
						Mout   <= ALU_CMP_OUT;
						CCR(2) <= ALU_CMP_CARRY;

					WHEN "10011" =>
						Mout   <= ALU_LDM_OUT;
						CCR(2) <= ALU_LDM_CARRY;

					WHEN OTHERS =>
						Mout <= (OTHERS => '0');
						CCR(2) <= '0';
				END CASE;
			END IF;
		END PROCESS;

		-- ZERO FLAG
		CCR(0) <= '1' WHEN (signed(Mout) = 0) ELSE '0';
		-- NEGATIVE FLAG
		CCR(1) <= '1' WHEN (signed(Mout) < 0) ELSE '0';

END a_OurALU;
