LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MIPS_Processor IS
	PORT (
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		
		Addrtest: IN STD_LOGIC_VECTOR(11 DOWNTO 0);

		DataOutTest : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END MIPS_Processor;

ARCHITECTURE a_MIPS_Processor OF MIPS_Processor IS

	COMPONENT PCount IS
		PORT (
			CLK : IN STD_LOGIC;
			RST : IN STD_LOGIC;
			NewValue : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Outdata  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT InstrCache IS
		PORT (
			Addr  : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    			Instruction  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT FetchDecode IS
		PORT (
			CLK : IN STD_LOGIC;
			RST : IN STD_LOGIC;
			NewValue : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			Outdata  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;

	SIGNAL PC : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PCout : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL INST : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL INSTBuf : STD_LOGIC_VECTOR(15 DOWNTO 0);

	BEGIN

		PC <= "00000000000000000000" & Addrtest;

		u0: PCount PORT MAP(CLK, RST, PC, PCout);
		u1: InstrCache PORT MAP(PCout(11 DOWNTO 0), INST);
		u2: FetchDecode PORT MAP(CLK, RST, INST, INSTBuf);
		

END a_MIPS_Processor;