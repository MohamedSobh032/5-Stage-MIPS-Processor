LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY PCount IS
	PORT (
		CLK      : IN  STD_LOGIC;
		RST      : IN  STD_LOGIC;
		ResetVal : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		NewValue : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Outdata  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END PCount;

ARCHITECTURE a_PCount OF PCount IS
	-- REGISTER --
    	SIGNAL PC : STD_LOGIC_VECTOR(31 DOWNTO 0);

	BEGIN
		PROCESS (CLK, RST)
		BEGIN
			IF (RST = '1') THEN
				PC <= ResetVal;
			ELSIF rising_edge(CLK) THEN
				PC <= NewValue;
			END IF;
		END PROCESS;	
		OutData <= PC;
END a_PCount;