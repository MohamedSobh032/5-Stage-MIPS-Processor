LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MIPS_Processor IS
	PORT (
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		INT : IN STD_LOGIC
	);
END MIPS_Processor;

ARCHITECTURE a_MIPS_Processor OF MIPS_Processor IS

	COMPONENT PCount IS
		PORT (
			CLK : IN STD_LOGIC;
			RST : IN STD_LOGIC;
			NewValue : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			Outdata  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT InstrCache IS
		PORT (
			Addr  : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    			Instruction  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT FetchDecode IS
		PORT (
			CLK : IN STD_LOGIC;
			RST : IN STD_LOGIC;
			NewValue : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			Outdata  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;

	BEGIN



END a_MIPS_Processor;