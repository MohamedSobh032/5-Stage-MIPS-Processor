LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY registerfile IS
	PORT (
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;

		-- decode stage
		Rsrc1 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Rsrc2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Rsrc1Data : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		Rsrc2Data : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);

		-- write back
		WE       : IN STD_LOGIC;
		Rdst     : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		RdstData : IN STD_LOGIC_VECTOR(31 DOWNTO 0);

	);
END registerfile;