LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY ControlUnit IS
	PORT (
		---------------- INSTRUCTION OPCODE ----------------
		INSTRUCTION : IN STD_LOGIC_VECTOR(4 DOWNTO 0);

		---------------- CONTROL SIGNALS ----------------
		-- WRITE BACK 1 		--> 0
		-- WRITE BACK 2 		--> 1
		-- Z/N F			--> 2
		-- C/OV F      		 	--> 3
		-- MemRead			--> 4
		-- MemWrite			--> 5
		-- FREE				--> 6
		-- PROTECT			--> 7
		-- IMMEDIATE			--> 8
		-- BRANCH			--> 9
		-- BRANCH ZERO 			--> 10
		-- SP DEC 			--> 11
		-- SP INC 		     	--> 12
		-- OUTPUT PORT   	     	--> 13
		-- INPUT PORT   	     	--> 14
		-- STORE                     	--> 15
		-- PUSH PC  	     		--> 16
		-- LENGTH EXT    	     	--> 17
		-- First Operand Dependency  	--> 18
		-- Second Operand Dependency 	--> 19
		-- PUSH CCR  			--> 20
		-- UPDATE PC USING MEMORY	--> 21
		-- POP CCR			--> 22
		CONTROL_SIGNALS : OUT STD_LOGIC_VECTOR(22 DOWNTO 0);

		---------------- ALU OPCODE ----------------
		-- NOT  --> 0001
		-- NEG  --> 0010
		-- INC  --> 0011
		-- DEC  --> 0100
		-- ADD  --> 0101
		-- ADDI --> 0101
		-- SUB  --> 0110
		-- SUBI --> 0110
		-- AND  --> 0111
		-- OR   --> 1000
		-- XOR  --> 1001
		-- CMP  --> 1010
		-- LDM  --> 1011
		-- LDD  --> 0101
		-- STD  --> 0101
		-- JZ   --> 1111
		ALU_OPCODE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE a_ControlUnit OF ControlUnit IS
	BEGIN
		---- ALU OPCODE SIGNAL SELECTION ----
		WITH INSTRUCTION SELECT
			ALU_OPCODE <=
				"0001" WHEN "00001", -- NOT
				"0010" WHEN "00010", -- NEG
				"0011" WHEN "00011", -- INC
				"0100" WHEN "00100", -- DEC
				"0101" WHEN "01001", -- ADD
				"0101" WHEN "01010", -- ADDI
				"0110" WHEN "01011", -- SUB
				"0110" WHEN "01100", -- SUBI
				"0111" WHEN "01101", -- AND
				"1000" WHEN "01110", -- OR
				"1001" WHEN "01111", -- XOR
				"0110" WHEN "10000", -- CMP
				"1011" WHEN "10011", -- LDM
				"0101" WHEN "10100", -- LDD
				"0101" WHEN "10101", -- STD
				"1111" WHEN "11000", -- JZ
				"0000" WHEN OTHERS;
		
		---- CONTROL SIGNAL SELECTION ----
		WITH INSTRUCTION SELECT
			CONTROL_SIGNALS <=
				"00000000000000000000000" WHEN "00000",	-- NOP
				"00001000000000000000101" WHEN "00001",	-- NOT
				"00001000000000000001101" WHEN "00010",	-- NEG
				"00001000000000000001101" WHEN "00011",	-- INC
				"00001000000000000001101" WHEN "00100",	-- DEC
				"00001000010000000000000" WHEN "00101",	-- OUT
				"00000000100000000000001" WHEN "00110",	-- IN
				"00001000000000000000001" WHEN "00111",	-- MOV
				"00001000000000000000011" WHEN "01000",	-- SWAP
				"00011000000000000001101" WHEN "01001",	-- ADD
				"00001000000000100001101" WHEN "01010",	-- ADDI
				"00011000000000000001101" WHEN "01011",	-- SUB
				"00001000000000100001101" WHEN "01100",	-- SUBI
				"00011000000000000000101" WHEN "01101",	-- AND
				"00011000000000000000101" WHEN "01110",	-- OR
				"00011000000000000000101" WHEN "01111",	-- XOR
				"00011000000000000000100" WHEN "10000",	-- CMP
				"00001000000100000100000" WHEN "10001",	-- PUSH
				"00000000001000000010001" WHEN "10010",	-- POP
				"00000100000000100000001" WHEN "10011",	-- LDM
				"00011000000000100010001" WHEN "10100",	-- LDD
				"00011001000000100100000" WHEN "10101",	-- STD
				"00000000000000010000000" WHEN "10110",	-- PROT
				"00000000000000001000000" WHEN "10111",	-- FREE
				"00001000000010000000100" WHEN "11000",	-- JZ
				"00001000000001000000000" WHEN "11001",	-- JMP
				"00001010000101000100000" WHEN "11010",	-- CALL
				"01000010001000000010000" WHEN "11011",	-- RET
				"01000010001000000010000" WHEN "11100",	-- RTI
				"00000010000100000100000" WHEN "11101", -- PUSH PC
				"00100000000100000100000" WHEN "11110", -- PUSH CCR
				"10000000001000000010000" WHEN "11111", -- POP THE CCR
				(OTHERS => '0') WHEN OTHERS;

END a_ControlUnit;
