LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY StackPointer IS
	PORT (
		CLK       : IN STD_LOGIC;
		RST       : IN STD_LOGIC;
		SP_INC    : IN STD_LOGIC;
		SP_DEC    : IN STD_LOGIC;
		SP_OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END StackPointer;

ARCHITECTURE a_StackPointer OF StackPointer IS
	-- REGISTER --
    	SIGNAL SP : STD_LOGIC_VECTOR(31 DOWNTO 0);

	-- LOGIC --
	SIGNAL SP_ADD_TWO : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SP_SUB_TWO : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SP_STAY    : STD_LOGIC_VECTOR(31 DOWNTO 0);

	-- OUTPUT SIGNAL --
	SIGNAL SP_TO_BE_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);

	BEGIN
		SP_ADD_TWO <= std_logic_vector(unsigned(SP) + 2);
		SP_SUB_TWO <= std_logic_vector(unsigned(SP) - 2);
		SP_STAY    <= SP;

		PROCESS (CLK, RST)
		BEGIN
			IF (RST = '1') THEN
				SP           <= x"FFFFFFFE";
				SP_TO_BE_OUT <= x"FFFFFFFE";
			ELSIF rising_edge(CLK) THEN

				IF (SP_INC = '1') THEN
					SP_TO_BE_OUT <= SP_ADD_TWO;
					SP           <= SP_ADD_TWO;
				END IF;

				IF (SP_DEC = '1') THEN
					SP_TO_BE_OUT <= SP_SUB_TWO;
					SP           <= SP_SUB_TWO;
				END IF;

			END IF;
		END PROCESS;
		SP_OUTPUT <= SP_TO_BE_OUT;
END a_StackPointer;

