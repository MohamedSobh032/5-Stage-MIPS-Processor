LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY PCount IS
	PORT (
		CLK      : IN  STD_LOGIC;
		RST      : IN  STD_LOGIC;
		INT      : IN  STD_LOGIC;
		EXCP     : IN  STD_LOGIC;
		PAUSE    : IN  STD_LOGIC;
		ResetVal : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		IntptVal : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		EXCPVal  : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		NewValue : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Outdata  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END PCount;

ARCHITECTURE a_PCount OF PCount IS
	-- REGISTER --
    	SIGNAL PC : STD_LOGIC_VECTOR(31 DOWNTO 0);

	BEGIN
		PROCESS (CLK, RST)
		BEGIN
			IF (RST = '1') THEN
				PC <= ResetVal;
			ELSIF (INT = '1') THEN
				PC <= IntptVal;
			ELSIF (EXCP = '1') THEN
				PC <= EXCPVal;
			ELSIF rising_edge(CLK) THEN
				IF (PAUSE = '0') THEN
					PC <= NewValue;
				END IF;
			END IF;
		END PROCESS;	
		OutData <= PC;
END a_PCount;