LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU_ldm IS
	PORT (
		Rsrc : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Rdst : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ALU_ldm;

ARCHITECTURE a_ALU_ldm OF ALU_ldm IS
	
	BEGIN
		Rdst <= Rsrc;

END a_ALU_ldm;