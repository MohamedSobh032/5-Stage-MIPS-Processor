LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU_mov IS
	PORT (
		Rsrc : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Rdst : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		Carry : OUT STD_LOGIC
	);
END ALU_mov;

ARCHITECTURE a_ALU_mov OF ALU_mov IS	
	BEGIN
		Rdst <= Rsrc;
		Carry <= '0';
END a_ALU_mov;
