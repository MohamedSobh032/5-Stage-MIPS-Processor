LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY StackPointer IS
	PORT (
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		NewValue : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Outdata  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END StackPointer;

ARCHITECTURE a_StackPointer OF StackPointer IS
    	SIGNAL SP : STD_LOGIC_VECTOR(31 DOWNTO 0);
	BEGIN
		PROCESS (CLK, RST)
		BEGIN
			IF (RST = '1') THEN
				SP <= (OTHERS => '1');
			ELSIF rising_edge(CLK) THEN
				SP <= NewValue;
			END IF;
		END PROCESS;	
		OutData <= SP;
END a_StackPointer;
