LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY JumpForwardUnit IS
	PORT (
		Rsrc_IN_E  : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Rdst_IN_WB : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		ZF_IN_WB   : IN STD_LOGIC;
		MR_IN_WB   : IN STD_LOGIC;
		ENABLE_BRANCHING : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE a_JumpForwardUnit OF JumpForwardUnit IS
	SIGNAL COMPARATOR : STD_LOGIC;
	BEGIN

		COMPARATOR <= '1' WHEN (Rsrc_IN_E = Rdst_IN_WB)
		ELSE          '0';
		ENABLE_BRANCHING <= COMPARATOR and ZF_IN_WB and MR_IN_WB;

END ARCHITECTURE;
