LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU_not IS
	PORT (
		Rsrc : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Rdst : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ALU_not;

ARCHITECTURE a_ALU_not OF ALU_not IS
	BEGIN
		Rdst <= not Rsrc;
END a_ALU_not;