LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DataForwardUnit IS
	PORT (
		Rsrc1Addr : IN STD_LOGIC_VECTOR(2 DOWNTO 0);

		Rdst1Addr_MEM   : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Rdst2Addr_MEM   : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		MEM_READ_IN_MEM : IN STD_LOGIC;
		SWAP_IN_MEM     : IN STD_LOGIC;

		Rdst1Addr_WB    : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Rdst2Addr_WB    : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		MEM_READ_IN_WB  : IN STD_LOGIC;
		SWAP_IN_WB      : IN STD_LOGIC
	);
END DataForwardUnit;


ARCHITECTURE a_DataForwardUnit OF DataForwardUnit IS

	BEGIN

		PROCESS (MEM_READ_IN_MEM, SWAP_IN_MEM, MEM_READ_IN_WB, SWAP_IN_WB)
		BEGIN
			IF (Rsrc1Addr = Rdst1Addr_MEM) THEN
				-- DATA FORWARD ALU-ALU
			ELSIF (Rsrc1Addr = Rdst2Addr_MEM) THEN
				-- DATA FORWARD ALU-ALU
				IF (SWAP_IN_MEM = '1') THEN

				END IF;
			END IF;
		END PROCESS;

END ARCHITECTURE;