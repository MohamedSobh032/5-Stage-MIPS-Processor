LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY OurALU IS
	PORT(
		CLK: IN STD_LOGIC;
		OPERATION: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		OP1, OP2: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		RESULT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		FLAGS: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END OurALU;

ARCHITECTURE a_OurALU OF OurALU IS

	SIGNAL S: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL F: STD_LOGIC_VECTOR(3 DOWNTO 0);

	BEGIN
		WITH OPERATION SELECT
			S <=
				NOT OP1 						     			   WHEN "0001", -- NOT
				STD_LOGIC_VECTOR(TO_SIGNED(0 - TO_INTEGER(SIGNED(OP1)), 32))	 		   WHEN "0010", -- NEG
				STD_LOGIC_VECTOR(TO_SIGNED(TO_INTEGER(SIGNED(OP1)) + 1, 32))			   WHEN "0011", -- INC
				STD_LOGIC_VECTOR(TO_SIGNED(TO_INTEGER(SIGNED(OP1)) - 1, 32)) 			   WHEN "0100", -- DEC
				STD_LOGIC_VECTOR(TO_SIGNED(TO_INTEGER(SIGNED(OP1)) + TO_INTEGER(SIGNED(OP2)), 32)) WHEN "0101", -- ADD
				STD_LOGIC_VECTOR(TO_SIGNED(TO_INTEGER(SIGNED(OP1)) - TO_INTEGER(SIGNED(OP2)), 32)) WHEN "0110", -- SUB
				OP1 AND OP2									   WHEN "0111", -- AND
				OP1 OR OP2									   WHEN "1000", -- OR
				OP1 XOR OP2									   WHEN "1001", -- XOR
				OP2										   WHEN "1011", -- LDM
				OP1										   WHEN OTHERS;

		F(3) <= '1' WHEN
				(OPERATION = "0010" AND '0' /= OP1(31) AND S(31) = OP1(31))
				OR (OPERATION = "0011" AND OP1(31) = '0' AND S(31) /= OP1(31))
				OR (OPERATION = "0100" AND OP1(31) /= '0' AND S(31) = '0')
				OR (OPERATION = "0101" AND OP1(31) = OP2(31) AND S(31) /= OP1(31))
				OR (OPERATION = "0110" AND OP1(31) /= OP2(31) AND S(31) = OP2(31))
		ELSE '0';

		F(2) <= '1' WHEN
			(OPERATION = "0010" AND 0 < TO_INTEGER(SIGNED(OP1)))
			OR (OPERATION = "0011" AND ((TO_INTEGER(SIGNED(S)) < TO_INTEGER(SIGNED(OP1))) OR (TO_INTEGER(SIGNED(S)) < 1)))
			OR (OPERATION = "0100" AND TO_INTEGER(SIGNED(OP1)) < 1)
			OR (OPERATION = "0101" AND ((TO_INTEGER(SIGNED(S)) < TO_INTEGER(SIGNED(OP1))) OR (TO_INTEGER(SIGNED(S)) < TO_INTEGER(SIGNED(OP2)))))
			OR (OPERATION = "0110" AND TO_INTEGER(SIGNED(OP1)) < TO_INTEGER(SIGNED(OP2)))
		ELSE '0';

		F(1) <= S(31);
		F(0) <= '1' WHEN S = X"00000000" ELSE '0';
		RESULT <= S;
		FLAGS <= F;
END a_OurALU;





