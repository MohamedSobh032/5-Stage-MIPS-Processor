LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY InReg IS
	PORT (
		Data_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		OutputPort : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END InReg;

ARCHITECTURE a_InReg OF InReg IS
	BEGIN
		OutputPort <= Data_IN;
END a_InReg;
