LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU_or IS
	PORT (
		Rsrc1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Rsrc2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Rdst  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ALU_or;

ARCHITECTURE a_ALU_or OF ALU_or IS
	BEGIN
		Rdst <= Rsrc1 or Rsrc2;
END a_ALU_or;